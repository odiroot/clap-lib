module clap

// String capacity for names that can be displayed to the user.
pub const name_size = 256
// String capacity for describing a path, like a parameter in a module
// hierarchy or path within a set of nested track groups.
pub const path_size = 1024
