module clap

pub type Id = u32

pub const invalid_id = Id(u32(C.CLAP_INVALID_ID))

