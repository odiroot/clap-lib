module clap

#flag -I @VMODROOT/include
#include "clap/clap.h"
